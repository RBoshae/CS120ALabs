`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:37:15 02/27/2017 
// Design Name: 
// Module Name:    timer_st 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module timer_st #( 
  parameter NBITS = 32  
)  
( 
   output wire timer ,  
   input wire  clk , 
   input wire  reset, 
   input [NBITS-1:0] cnt_ini ,   
   input [NBITS-1:0] cnt_rst   
 
);  

 
wire [NBITS-1:0] q ;    
wire [NBITS-1:0] qnext ;  
 
// Compute the next value  
 
adder #( .NBITS(NBITS ) )  
      c1 (.q(q),  
   .cnt_ini(cnt_ini),  
   .cnt_rst(cnt_rst),  
   .nextq(qnext),  
   .tick(timer) );  
 
// Save the next state  
flopr #( .NBITS(NBITS ) )  
      c2 (.clk(clk),  
  .reset(reset),  
   .cnt_ini(cnt_ini),  
   .nextq(qnext),  
   .q(q) ); 
 
endmodule 
