// Verilog test fixture created from schematic C:\Users\rwbos\Documents\GitHub\CS120ALabs\Lab5\datapath_components_adders_parta\four_bit_ripple_carry_adder.sch - Fri Feb 24 16:57:08 2017

`timescale 1ns / 1ps

module four_bit_ripple_carry_adder_four_bit_ripple_carry_adder_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   four_bit_ripple_carry_adder UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
