// Verilog test fixture created from schematic C:\Users\KongK\Documents\GitHub\CS120ALabs\Lab4\rising_edge_detector\rising_edge_detector_sm.sch - Mon Feb 13 15:56:32 2017

`timescale 1ns / 1ps

module rising_edge_detector_sm_rising_edge_detector_sm_sch_tb();

// Inputs
	reg signal;
	reg clk;
	
// Output
	wire outedge;
	
// Bidirs

// Instantiate the UUT
   rising_edge_detector_sm UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
